module miniproject(
);

endmodule